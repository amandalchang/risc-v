// given op, creates immSrc to control the immediate extender
/*
immSrc  | immExt
  00    |
  01    |
  10    |
  11    |


*/

module instruction_decoder(
    input logic clk,
    input [6:0] op,
    output [1:0] immsrc
);

endmodule