// Control Unit
// given the op code, funct3, and funct7, outputs control signals to the rest of the processor

`include "alu_decoder.sv"
`include "instr_decoder.sv"


module control(
    output logic    pc_write,
    output logic    adr_src,
    output logic    mem_write,
    output logic    ir_write,
    input logic     clk,
    input logic     [31:0] instr,
    input logic     zero,
    input logic     carry,
    input logic     negative,
    input logic     overflow,
    output logic    [1:0] result_src,
    output logic    [3:0] alu_control,
    output logic    [1:0] alu_src_b,
    output logic    [1:0] alu_src_a,
    output logic    [2:0] imm_src,
    output logic    reg_write
);

    logic [6:0] opcode;
    logic [2:0] funct3;
    logic [6:0] funct7;

    assign opcode = instr[6:0];
    assign funct3 = instr[14:12];
    assign funct7 = instr[31:25];

    logic pc_update = 1'b0;
    logic branch = 1'b0;
    logic [1:0] alu_op;
    // State variables
    localparam [2:0] FETCH = 3'b000;
    localparam [2:0] DECODE = 3'b001;
    localparam [2:0] EXECUTE = 3'b010;
    localparam [2:0] MEMORY = 3'b011;
    localparam [2:0] WRITE_BACK = 3'b100;

    // opcodes
    localparam [6:0] LOAD = 7'b0000011;
    localparam [6:0] STORE = 7'b0100011;
    localparam [6:0] EXECUTE_R = 7'b0110011;
    localparam [6:0] EXECUTE_I = 7'b0010011;
    localparam [6:0] JAL = 7'b1101111;
    localparam [6:0] JALR = 7'b1100111;
    localparam [6:0] BRANCH = 7'b1100011;
    localparam [6:0] EXECUTE_LUI = 7'b0110111;
    localparam [6:0] EXECUTE_AUIPC = 7'b0010111;
    
    // alu_src_a and alu_src_b localparams
    localparam [1:0] A_SELECT_PC = 2'b00;
    localparam [1:0] A_SELECT_OLD_PC = 2'b01;
    localparam [1:0] A_SELECT_RD1 = 2'b10;

    localparam [1:0] B_SELECT_RD2 = 2'b00;
    localparam [1:0] B_SELECT_IMM_EXT = 2'b01;
    localparam [1:0] B_SELECT_4 = 2'b10;

    // alu_op localparams
    localparam [1:0] ADD = 2'b00;
    localparam [1:0] SUB = 2'b01;
    localparam [1:0] FUNCT3_DEPEND = 2'b10;
    localparam [1:0] PASS = 2'b11;


    // Declare state variables
    logic [2:0] current_state = FETCH;

    // Thus, the N (Negative) flag is connected to the most significant bit of the ALU output, Result31. 
// The Z (Zero) flag is asserted when all of the bits of Result are 0, as detected by the N-bit NOR gate in Figure 5.17. 
// The C (Carry out) flag is asserted when the adder produces a carry out
//          and the ALU is performing addition or subtraction (indicated by ALUControl1 = 0).
// logic zero;
// logic carry;
// logic negative;
// WHEN THESE 3 THINGS ARE TRUE
// (1) the ALU is performing addition or subtraction (ALUControl1 = 0)
// (2) A and Sum have opposite signs, as detected by the XOR gate
// (3) overflow is possible. That is, as detected by the XNOR gate, either A and B have the same negative 
//          and the adder is performing addition (ALUControl0 = 0) or A and B have opposite signs 
//          and the adder is performing subtraction (ALUControl0 = 1). 
    


    always_ff @(posedge clk) begin
        if (current_state == WRITE_BACK) begin
            current_state <= FETCH;
        end else begin
            current_state <= current_state + 1'b1;
        end
    end

    always_comb begin
        pc_update = 1'b0;
        branch = 1'b0;
        reg_write = 1'b0;
        ir_write = 1'b0;
        mem_write = 1'b0;
        // if it's time to increment
        case (current_state) // increment based on state
            FETCH: begin
                // reset enables
                reg_write = 1'b0;
                mem_write = 1'b0;
                branch = 1'b0;
                // state logic
                adr_src = 1'b0;
                ir_write = 1'b1;
                alu_src_a = A_SELECT_PC; // pc
                alu_src_b = B_SELECT_4; // 4
                alu_op = ADD; // ADD
                result_src = 2'b10; // from ALUResult
                pc_update = 1'b1; // prep for jump/branch
            end
            DECODE: begin
                // reset enables
                ir_write = 1'b1;
                pc_update = 1'b0;
                // state logic
                alu_src_a = A_SELECT_OLD_PC;
                alu_src_b = B_SELECT_IMM_EXT;
                alu_op = ADD;
            end
            EXECUTE: begin
                case(opcode)
                    LOAD, STORE: begin
                        alu_src_a = A_SELECT_RD1;
                        alu_src_b = B_SELECT_IMM_EXT;
                        alu_op = ADD;
                        adr_src = 1'b1;
                    end
                    EXECUTE_R: begin
                        // state logic
                        alu_src_a = A_SELECT_RD1;
                        alu_src_b = B_SELECT_RD2;
                        alu_op = FUNCT3_DEPEND;
                    end
                    EXECUTE_I: begin
                        // state logic
                        alu_src_a = A_SELECT_RD1;
                        alu_src_b = B_SELECT_IMM_EXT;
                        alu_op = FUNCT3_DEPEND;
                    end
                    JAL: begin
                        // state logic
                        alu_src_a = A_SELECT_OLD_PC;
                        alu_src_b = B_SELECT_4;
                        alu_op = ADD;
                        result_src = 2'b00;
                        pc_update = 1'b1;
                    end
                    JALR: begin
                        alu_src_a = A_SELECT_OLD_PC;
                        alu_src_b = B_SELECT_4;
                        alu_op = ADD;
                        result_src = 2'b10;
                        reg_write = 1'b1;
                    end
                    BRANCH: begin
                        // state logic
                        alu_src_a = A_SELECT_RD1;
                        alu_src_b = B_SELECT_RD2;
                        alu_op = SUB;
                        result_src = 2'b00;
                        branch = 1'b1;
                    end
                    EXECUTE_LUI: begin
                        alu_src_b = B_SELECT_IMM_EXT;
                        alu_op = PASS;
                        result_src = 2'b10;
                        reg_write = 1'b1;
                    end
                    EXECUTE_AUIPC: begin
                        alu_src_b = B_SELECT_IMM_EXT;
                        alu_op = ADD;
                        result_src = 2'b10;
                        reg_write = 1'b1;
                    end
                    default: begin
                        // Do nothing
                    end
                endcase
            end
            MEMORY: begin
                case(opcode)
                    LOAD: begin
                        result_src = 2'b00;
                        adr_src = 1'b1;
                    end
                    STORE: begin
                        result_src = 2'b00;
                        adr_src = 1'b1;
                        mem_write = 1'b1;
                    end
                    EXECUTE_R, EXECUTE_I, JAL: begin // ALUWB
                        result_src = 2'b00;
                        reg_write = 1'b1;
                    end
                    JALR: begin
                        alu_src_a = A_SELECT_RD1;
                        alu_src_b = B_SELECT_IMM_EXT;
                        alu_op = ADD;
                        result_src = 2'b10;
                        pc_update = 1'b1;
                    end
                    STORE: begin
                        result_src = 2'b00;
                        adr_src = 1'b1;
                        mem_write = 1'b1;
                    end
                    default: begin
                        // Do nothing
                    end
                endcase
            end
            WRITE_BACK: begin
                if (opcode == LOAD) begin
                    result_src = 2'b01;
                    reg_write = 1'b1;
                    adr_src = 1'b0;
                end
            end
        endcase
    end

    always_comb begin
        pc_write = pc_update;
        if (branch) begin
            case (funct3)
                3'b000: pc_write = zero; // BEQ
                3'b001: pc_write = !zero; // BNEQ
                3'b100: pc_write = negative; // BLT
                3'b101: pc_write = !negative; // BGE
                3'b110: pc_write = carry; // BLTU
                3'b111: pc_write = !carry; // BGEU
            endcase
        end
    end

    ALU_decoder ALU_decoder (
        .clk            (clk), 
        .funct3         (funct3),
        .op_5           (opcode[5]),
        .funct7_5       (funct7[5]),
        .alu_op         (alu_op),
        .alu_control    (alu_control)

    );

    instruction_decoder instruction_decoder (
        .clk            (clk), 
        .op             (opcode),
        .imm_src        (imm_src)
    );

endmodule